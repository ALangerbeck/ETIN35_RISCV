library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity stage_ex is
    generic(DATA_WIDTH: integer := 32);

    port(
        Data  : inout std_logic
    );
end stage_ex;

architecture behavioral of stage_ex is


begin



end behavioral;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity stage_id is
    generic(DATA_WIDTH: integer := 32);

    port(
        
    );
end stage_id;

architecture behavioral of stage_id is


begin



end behavioral;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;

entity stage_wb is
    port(
        ALU_result : in std_logic_vector(DATA_WIDTH-1 downto 0)
        
    );
end stage_wb;

architecture behavioral of stage_wb is


begin



end behavioral;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity stage_if is
    generic(DATA_WIDTH: integer := 32);

    port(
        
    );
end stage_if;

architecture behavioral of stage_if is


begin



end behavioral;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;
use STD.textio.all;

entity risc_v_tb is
end entity;


architecture structural of  risc_v_tb is


	--Signal Declaration

	--Component declaration

	
begin
  

end structural;
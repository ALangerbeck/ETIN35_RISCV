library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity stage_mem is
    generic(DATA_WIDTH: integer := 32);

    port(
        
    );
end stage_mem;

architecture behavioral of stage_mem is


begin



end behavioral;